module BROM(
    input ck;
    input [DATA_WIDTH:0] addr;
    input [DATA_WIDTH:0] din;
    input wen;
    output [DATA_WIDTH:0] dout;
);

endmodule // BROM